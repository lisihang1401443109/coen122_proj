module datapath_test (

);

    
endmodule